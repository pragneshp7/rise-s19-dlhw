import FIFO::*;

(* synthesize *)
module mkTop ();

    rule finish_sim;
        $display("Hello Priyal12");
        $finish;
    endrule
endmodule
